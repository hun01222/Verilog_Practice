module new;
  initial begin
    $display("hello world !");
  end
endmodule