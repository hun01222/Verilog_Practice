module t_flip_flop_structural_module(t, clk, q, q_bar);
  input t;
  input clk;

  output q, q_bar;
  reg q, q_bar;


endmodule