//This is for the D latch module.

module d_latch_gatelevel_module (d, en, q, q_bar);
	input d;
	input en; //enable

	output q, q_bar;
	
	wire not_1_output;
	wire and_1_output, and_2_output;
	wire or_1_output, or_2_output;
	
	//Fill this out.
	
endmodule
