//This is for the 4:2 priority encoder module.

module four_to_two_priority_encoder_gatelevel_module (a, b, c, d, out0, out1);
	input a, b, c, d;

	output out0, out1;
	
	//Fill this out

endmodule
