//This is for the D latch module.

module d_latch_sturctural_module (d, en, q, q_bar);
	input d;
	input en; //enable

	output q, q_bar;
	
	wire not_1_output;
	
	//Fill this out.
	
endmodule

