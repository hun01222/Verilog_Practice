module instructionMemory_P1
    #(parameter Width = 32)
(
    input  [Width-1:0] address,
    output [Width-1:0] instruction
);
    reg [9:0] cutAddress;
    reg [Width-1:0] mem[0:1023];

    initial begin
        //lw
        mem[ 0] = 32'h0078783; //lw  mem[x15]->x15 000000000000 01111 000 01111 0000011
        mem[ 4] = 32'h0080803; //lw  mem[x16]->x16 000000000000 10000 000 10000 0000011
        mem[ 8] = 32'h0088883; //lw  mem[x17]->x17 000000000000 10001 000 10001 0000011
        mem[12] = 32'h0090903; //lw  mem[x18]->x18 000000000000 10010 000 10010 0000011
        mem[16] = 32'h0098983; //lw  mem[x19]->x19 000000000000 10011 000 10011 0000011
        mem[20] = 32'h00A0A03; //lw  mem[x20]->x20 000000000000 10100 000 10100 0000011
        mem[24] = 32'h00A8A83; //lw  mem[x21]->x21 000000000000 10101 000 10101 0000011
        mem[28] = 32'h00B0B03; //lw  mem[x22]->x22 000000000000 10110 000 10110 0000011
        mem[32] = 32'h00B8B83; //lw  mem[x23]->x23 000000000000 10111 000 10111 0000011
        mem[36] = 32'h00C0C03; //lw  mem[x24]->x24 000000000000 11000 000 11000 0000011
        mem[40] = 32'h00C8C83; //lw  mem[x25]->x25 000000000000 11001 000 11001 0000011
        mem[44] = 32'h00D0D03; //lw  mem[x26]->x26 000000000000 11010 000 11010 0000011
        
        //R-type
        mem[48] = 32'h40FC1DB3; //mul x27,x15,x24 0100000 01111 11000 001 11011 0110011
        mem[52] = 32'h410C95B3; //mul x11,x16,x25 0100000 10000 11001 001 01011 0110011
        mem[56] = 32'h00BD8DB3; //add x27,x11,x27 0000000 01011 11011 000 11011 0110011
        mem[60] = 32'h411D15B3; //mul x11,x17,x26 0100000 10001 11010 001 01011 0110011
        mem[64] = 32'h00BD8DB3; //add x27,x11,x27 0000000 01011 11011 000 11011 0110011

        mem[68] = 32'h412C1E33; //mul x28,x18,x24 0100000 10010 11000 001 11100 0110011
        mem[72] = 32'h413C95B3; //mul x11,x19,x25 0100000 10011 11001 001 01011 0110011
        mem[76] = 32'h00BE0E33; //add x28,x11,x28 0000000 01011 11100 000 11100 0110011
        mem[80] = 32'h414D15B3; //mul x11,x20,x26 0100000 10100 11010 001 01011 0110011
        mem[84] = 32'h00BE0E33; //add x28,x11,x28 0000000 01011 11100 000 11100 0110011

        mem[88] = 32'h415C1EB3; //mul x29,x21,x24 0100000 10101 11000 001 11101 0110011
        mem[92] = 32'h416C95B3; //mul x11,x22,x25 0100000 10110 11001 001 01011 0110011
        mem[96] = 32'h00BE8EB3; //add x29,x11,x29 0000000 01011 11101 000 11101 0110011
        mem[100] = 32'h417D15B3; //mul x11,x23,x26 0100000 10111 11010 001 01011 0110011
        mem[104] = 32'h00BE8EB3; //add x29,x11,x29 0000000 01011 11101 000 11101 0110011
        
        //store
        mem[108] = 32'h01B60007; //sw x27->mem[x12] 0000000 11011 01100 000 00000 0000111
        mem[112] = 32'h01C68007; //sw x28->mem[x13] 0000000 11100 01101 000 00000 0000111
        mem[116] = 32'h01D70007; //sw x29->mem[x14] 0000000 11101 01110 000 00000 0000111
    end
    assign instruction = mem[address];
endmodule
